`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// National University of Singapore
// Department of Electrical and Computer Engineering
// EE2026 Digital Design
// AY1819 Semester 1
// Project: Voice Scope
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////
// Menu
// hide elements(basic feature)
// circle improvement - layers
// ///////////////////////////
module Voice_Scope_TOP(
    input CLK, btnL, btnR, btnU, btnD, btnC,
    input [2:0] color_set,
    input [15:0] sw,
    input  J_MIC3_Pin3,   // PmodMIC3 audio input data (serial)
    output J_MIC3_Pin1,   // PmodMIC3 chip select, 20kHz sampling clock
    output J_MIC3_Pin4,   // PmodMIC3 serial clock (generated by module VoiceCapturer.v)
   
    output [3:0] VGA_RED,    // RGB outputs to VGA connector (4 bits per channel gives 4096 possible colors)
    output [3:0] VGA_GREEN,
    output [3:0] VGA_BLUE,
    output VGA_VS,          // horizontal & vertical sync outputs to VGA connector
    output VGA_HS,
    output [11:0] led,
    output [3:0] an,
    output [6:0] seg
    );
       
   
      
       
//-----------------------------------------------------------------------------
//                  STUDENT A - MIC
//-----------------------------------------------------------------------------
// Please create a clock divider module to generate a 20kHz clock signal. 
// Instantiate it below
    wire clk_20k;
    wire slow_clock;
    wire slower_clock;
    wire [11:0]gen_wave;
    clk_div a (CLK,clk_20k,slow_clock,slower_clock);
// Please instantiate the voice capturer module below
    Voice_Capturer b (CLK,clk_20k,J_MIC3_Pin3,J_MIC3_Pin1,J_MIC3_Pin4,gen_wave);

//-----------------------------------------------------------------------------
//                  STUDENT B - VGA
//-----------------------------------------------------------------------------
    wire [11:0] VGA_HORZ_COORD;
    wire [11:0] VGA_VERT_COORD; 
    wire [3:0] VGA_Red_waveform;
    wire [3:0] VGA_Green_waveform;
    wire [3:0] VGA_Blue_waveform;
    wire [9:0] wave_sample; 
    wire [9:0] test_wave_sample; 
    wire [3:0] VGA_Red_grid;
    wire [3:0] VGA_Green_grid;
    wire [3:0] VGA_Blue_grid;
    wire [3:0] VGA_Red_out;
    wire [3:0] VGA_Green_out;
    wire [3:0] VGA_Blue_out;
    wire [3:0] VGA_Red_Pong;
    wire [3:0] VGA_Green_Pong;
    wire [3:0] VGA_Blue_Pong;
    wire [3:0] VGA_Red_Intro;
    wire [3:0] VGA_Green_Intro;
    wire [3:0] VGA_Blue_Intro;
    wire [3:0] red_menu;
    wire [3:0] green_menu;
    wire [3:0] blue_menu;
    wire [3:0] red_pong;
    wire [3:0] green_pong;
    wire [3:0] blue_pong;    
    wire [3:0] red_bar;
    wire [3:0] green_bar;
    wire [3:0] blue_bar;
    wire [0:11] bg;
    wire [0:11] grid;
    wire [0:11] waveform;
    wire [0:11] tick;
    wire [0:11] axis;
    wire [3:0] lvl;
    wire up,down,center,left,right;
    wire [1:0]STATE;
    wire MAIN_MENU;
    wire [1:0]SIDE_MENU_GRAPH;
    wire SIDE_MENU_PONG;
    wire [1:0]GRAPH;
    wire PONG;
    wire [1:0]COLOR;
    wire wave_cond1,wave_cond2;
    wire menu_bg,color_box;
    
    wire [3:0] VGA_Red_waveform1;
    wire [3:0] VGA_Red_waveform2;
    wire [3:0] VGA_Red_waveform3;
    wire [3:0] VGA_Red_waveform4;
    wire [3:0] VGA_Red_waveform5;
    wire [3:0] VGA_Red_waveform6;
    wire [3:0] VGA_Red_waveform7;
    wire [3:0] VGA_Red_waveform8;
    wire [3:0] VGA_Red_waveform9;
    wire [3:0] VGA_Red_waveform10;
    wire [3:0] VGA_Red_waveform11;
    wire [3:0] VGA_Red_waveform12;
    wire [3:0] VGA_Red_waveform13;
    wire [3:0] VGA_Red_waveform14;
    wire [3:0] VGA_Red_waveform15;
    
    wire [3:0] VGA_Green_waveform1;
    wire [3:0] VGA_Green_waveform2;
    wire [3:0] VGA_Green_waveform3;
    wire [3:0] VGA_Green_waveform4;
    wire [3:0] VGA_Green_waveform5;
    wire [3:0] VGA_Green_waveform6;
    wire [3:0] VGA_Green_waveform7;
    wire [3:0] VGA_Green_waveform8;
    wire [3:0] VGA_Green_waveform9;
    wire [3:0] VGA_Green_waveform10;
    wire [3:0] VGA_Green_waveform11;
    wire [3:0] VGA_Green_waveform12;
    wire [3:0] VGA_Green_waveform13;
    wire [3:0] VGA_Green_waveform14;
    wire [3:0] VGA_Green_waveform15;
    
    wire [3:0] VGA_Blue_waveform1;
    wire [3:0] VGA_Blue_waveform2;
    wire [3:0] VGA_Blue_waveform3;
    wire [3:0] VGA_Blue_waveform4;
    wire [3:0] VGA_Blue_waveform5;
    wire [3:0] VGA_Blue_waveform6;
    wire [3:0] VGA_Blue_waveform7;
    wire [3:0] VGA_Blue_waveform8;
    wire [3:0] VGA_Blue_waveform9;
    wire [3:0] VGA_Blue_waveform10;
    wire [3:0] VGA_Blue_waveform11;
    wire [3:0] VGA_Blue_waveform12;
    wire [3:0] VGA_Blue_waveform13;
    wire [3:0] VGA_Blue_waveform14;
    wire [3:0] VGA_Blue_waveform15;

    wire [3:0] VGA_Red_grid1;
    wire [3:0] VGA_Red_grid2;
    wire [3:0] VGA_Red_grid3;
    wire [3:0] VGA_Red_grid4;
    wire [3:0] VGA_Red_grid5;
    wire [3:0] VGA_Red_grid6;
    wire [3:0] VGA_Red_grid7;
    wire [3:0] VGA_Red_grid8;
    wire [3:0] VGA_Red_grid9;
    wire [3:0] VGA_Red_grid10;
    wire [3:0] VGA_Red_grid11;
    wire [3:0] VGA_Red_grid12;
    wire [3:0] VGA_Red_grid13;
    wire [3:0] VGA_Red_grid14;
    wire [3:0] VGA_Red_grid15;
    
    wire [3:0] VGA_Green_grid1;
    wire [3:0] VGA_Green_grid2;
    wire [3:0] VGA_Green_grid3;
    wire [3:0] VGA_Green_grid4;
    wire [3:0] VGA_Green_grid5;
    wire [3:0] VGA_Green_grid6;
    wire [3:0] VGA_Green_grid7;
    wire [3:0] VGA_Green_grid8;
    wire [3:0] VGA_Green_grid9;
    wire [3:0] VGA_Green_grid10;
    wire [3:0] VGA_Green_grid11;
    wire [3:0] VGA_Green_grid12;
    wire [3:0] VGA_Green_grid13;
    wire [3:0] VGA_Green_grid14;
    wire [3:0] VGA_Green_grid15;
    
    wire [3:0] VGA_Blue_grid1;
    wire [3:0] VGA_Blue_grid2;
    wire [3:0] VGA_Blue_grid3;
    wire [3:0] VGA_Blue_grid4;
    wire [3:0] VGA_Blue_grid5;
    wire [3:0] VGA_Blue_grid6;
    wire [3:0] VGA_Blue_grid7;
    wire [3:0] VGA_Blue_grid8;
    wire [3:0] VGA_Blue_grid9;
    wire [3:0] VGA_Blue_grid10;
    wire [3:0] VGA_Blue_grid11;
    wire [3:0] VGA_Blue_grid12;
    wire [3:0] VGA_Blue_grid13;
    wire [3:0] VGA_Blue_grid14;
    wire [3:0] VGA_Blue_grid15;
    
    reg [3:0]graph_out_red;
    reg [3:0]graph_out_green;
    reg [3:0]graph_out_blue;
    assign VGA_Red_out = (STATE == 0) ? VGA_Red_Intro : (STATE == 1) ? graph_out_red|red_menu  : (STATE == 2) ? (red_pong|VGA_Red_Pong) : 0;
    assign VGA_Green_out = (STATE == 0) ?VGA_Green_Intro: (STATE == 1) ? graph_out_green|green_menu : (STATE == 2) ? (green_pong | VGA_Green_Pong) : 0;
    assign VGA_Blue_out = (STATE == 0) ? VGA_Blue_Intro: (STATE == 1) ? graph_out_blue|blue_menu: (STATE == 2)  ? (blue_pong | VGA_Blue_Pong) : 0;
    
    wire line_graph2 = (VGA_HORZ_COORD % 10 == 0);
    wire VGA_CLOCK;
    wire [4:0]GRAPH_STATE;
    wire zoom;
    wire [1:0]bar_size;
    
    
    always @ (posedge VGA_CLOCK)begin
        
        case(GRAPH_STATE)
            0:
            begin
                graph_out_red <= VGA_Red_grid | VGA_Red_waveform ;
                graph_out_green <=  VGA_Green_grid | VGA_Green_waveform ;
                graph_out_blue <= VGA_Blue_grid | VGA_Blue_waveform ;
            end
            1:
            begin
                graph_out_red <= VGA_Red_grid | VGA_Red_waveform | VGA_Red_grid9;
                graph_out_green <=  VGA_Green_grid | VGA_Green_waveform | VGA_Green_grid9;
                graph_out_blue <= VGA_Blue_grid | VGA_Blue_waveform | VGA_Blue_grid9;                
            end
            2:
            begin
                graph_out_red <= VGA_Red_waveform | VGA_Red_grid7;
                graph_out_green <= VGA_Green_waveform | VGA_Green_grid7;
                graph_out_blue <= VGA_Blue_waveform | VGA_Blue_grid7; 
            end
            3:
            begin
                graph_out_red <= VGA_Red_waveform8 | VGA_Red_grid8;
                graph_out_green <= VGA_Green_waveform8 | VGA_Green_grid8;
                graph_out_blue <= VGA_Blue_waveform8 | VGA_Blue_grid8;
            end
            4:
            begin
                graph_out_red <= red_bar;
                graph_out_green <= green_bar;
                graph_out_blue <= blue_bar;
            end
            5:
            begin
                graph_out_red <= red_bar;
                graph_out_green <= green_bar;
                graph_out_blue <= blue_bar;
            end
            6:
            begin
                graph_out_red <=  VGA_Red_grid4;
                graph_out_green <=  VGA_Green_grid4;
                graph_out_blue <=  VGA_Blue_grid4;
            end
            7:
            begin
                graph_out_red <= VGA_Red_grid1;
                graph_out_green <= VGA_Green_grid1;
                graph_out_blue <= VGA_Blue_grid1;
            end
            8:
            begin
                graph_out_red <= VGA_Red_grid2;
                graph_out_green <= VGA_Green_grid2;
                graph_out_blue <= VGA_Blue_grid2;
            end
            9:
            begin
                graph_out_red <= VGA_Red_waveform10 | VGA_Red_grid10;
                graph_out_green <= VGA_Green_waveform10 | VGA_Green_grid10;
                graph_out_blue <= VGA_Blue_waveform10 | VGA_Blue_grid10;
            end
            10:
            begin
                graph_out_red <= VGA_Red_waveform11 | VGA_Red_grid11;
                graph_out_green <= VGA_Green_waveform11 | VGA_Green_grid11;
                graph_out_blue <= VGA_Blue_waveform11 | VGA_Blue_grid11;
            end
            11:
            begin
                graph_out_red <= VGA_Red_waveform12 | VGA_Red_grid12;
                graph_out_green <= VGA_Green_waveform12 | VGA_Green_grid12;
                graph_out_blue <= VGA_Blue_waveform12 | VGA_Blue_grid12;
            end
            12:
            begin
                graph_out_red <= VGA_Red_waveform13 | VGA_Red_grid13;
                graph_out_green <= VGA_Green_waveform13 | VGA_Green_grid13;
                graph_out_blue <= VGA_Blue_waveform13 | VGA_Blue_grid13;
            end
            13:
            begin
                graph_out_red <= VGA_Red_waveform6 | VGA_Red_grid6;
                graph_out_green <= VGA_Green_waveform6 | VGA_Green_grid6;
                graph_out_blue <= VGA_Blue_waveform6 | VGA_Blue_grid6;
            end
            14:
            begin
                graph_out_red <= VGA_Red_waveform15 | VGA_Red_grid15;
                graph_out_green <= VGA_Green_waveform15 | VGA_Green_grid15;
                graph_out_blue <= VGA_Blue_waveform15 | VGA_Blue_grid15;
            end
        endcase
    end
    wire [0:11] input_color;
    assign wave_sample = sw[0] ? test_wave_sample : gen_wave >> 2;
    TestWave_Gen c (clk_20k,test_wave_sample);
    Draw_Waveform d(sw[10],zoom,waveform,clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform,VGA_Green_waveform,VGA_Blue_waveform,wave_cond1,wave_cond2);
    Draw_Background e(sw[10:7],SIDE_MENU_GRAPH,menu_bg,color_box,wave_cond1,axis,bg,grid,tick,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid,VGA_Green_grid,VGA_Blue_grid);
    Draw_Pong f (SIDE_MENU_PONG,menu_bg,STATE,lvl,slow_clock,sw[15],sw[3],sw[2],sw[14],sw[4],VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_Pong,VGA_Green_Pong,VGA_Blue_Pong);
    VGA_DISPLAY g(CLK,VGA_Red_out,VGA_Green_out,VGA_Blue_out,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_RED,VGA_GREEN,VGA_BLUE,VGA_VS,VGA_HS,VGA_CLOCK);
    color_select h(center,sw[13:11],input_color,SIDE_MENU_GRAPH,slow_clock,left,right,bg,grid,waveform,tick,axis);
    introduction i(MAIN_MENU,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_Intro,VGA_Green_Intro,VGA_Blue_Intro);
    menu_graph j(GRAPH_STATE,left,right,SIDE_MENU_GRAPH,GRAPH,COLOR,slow_clock,VGA_HORZ_COORD,VGA_VERT_COORD,red_menu,green_menu,blue_menu,menu_bg,color_box,input_color);
    menu_pong k(menu_bg,SIDE_MENU_PONG,PONG,VGA_HORZ_COORD,VGA_VERT_COORD,red_pong,green_pong,blue_pong);
    menu_logic l(up,down,center,slow_clock,STATE,MAIN_MENU,SIDE_MENU_GRAPH,SIDE_MENU_PONG,GRAPH,PONG,COLOR,GRAPH_STATE,zoom,bar_size);
    bar_graph m(bar_size,grid,clk_20k,wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,red_bar,green_bar,blue_bar);
    vert_zoom1b o(wave_cond1,slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid7,VGA_Green_grid7,VGA_Blue_grid7);
    full1 p(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform15,VGA_Green_waveform15,VGA_Blue_waveform15);
    full2 q(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], lvl, VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid15,VGA_Green_grid15,VGA_Blue_grid15);
    full3 p1(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform6,VGA_Green_waveform6,VGA_Blue_waveform6);
    full4 q2(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], lvl, VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid6,VGA_Green_grid6,VGA_Blue_grid6);
    line_graph1 e1(slower_clock,axis,bg,grid,tick,clk_20k,wave_cond2,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid6,VGA_Green_grid1,VGA_Blue_grid1);
    line_graph2 e2(slower_clock,axis,bg,grid,tick,clk_20k,wave_cond2,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid2,VGA_Green_grid2,VGA_Blue_grid2);
    
    vert_zoom2a d8(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform8,VGA_Green_waveform8,VGA_Blue_waveform8);
    vert_zoom2b e8(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid8,VGA_Green_grid8,VGA_Blue_grid8);
    
    volume_indicate e9(menu_bg,color_box,SIDE_MENU_GRAPH,slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid9,VGA_Green_grid9,VGA_Blue_grid9);
    
    slow_waveform1 d10(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform10,VGA_Green_waveform10,VGA_Blue_waveform10);
    slow_background1 e10(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid10,VGA_Green_grid10,VGA_Blue_grid10);
     
    slow_waveform2 d11(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform11,VGA_Green_waveform11,VGA_Blue_waveform11);
    slow_background2 e11(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid11,VGA_Green_grid11,VGA_Blue_grid11);

    display1 d12(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform12,VGA_Green_waveform12,VGA_Blue_waveform12);
    display2 e12(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid12,VGA_Green_grid12,VGA_Blue_grid12);
        
    display1 d13(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform13,VGA_Green_waveform13,VGA_Blue_waveform13);
    display3 e13(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid13,VGA_Green_grid13,VGA_Blue_grid13);
     
    horiz_display1 d14(bg,waveform, clk_20k,sw[1],wave_sample,VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_waveform14,VGA_Green_waveform14,VGA_Blue_waveform14);
    horiz_display2 e14(slower_clock,axis,bg,grid,tick,clk_20k,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid14,VGA_Green_grid14,VGA_Blue_grid14);

    draw_circle e3(axis,bg,grid,tick,clk_20k,lvl,wave_sample,sw[1], VGA_HORZ_COORD,VGA_VERT_COORD,VGA_Red_grid4,VGA_Green_grid4,VGA_Blue_grid4);

    debounce t(slow_clock,btnL,left);
    debounce u(slow_clock,btnR,right);
    debounce v(slow_clock,btnU,up);
    debounce w(slow_clock,btnD,down);
    debounce x(slow_clock,btnC,center);
    vol_indi y (wave_sample,clk_20k,led,lvl);
    sev_seg z(lvl,clk_20k,an,seg);
endmodule
